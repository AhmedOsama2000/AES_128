package aes_uvm_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	// Include UVM_CLASSES
	`include "Sequence_item.sv"
	`include "Sequence.sv"
	`include "Sequencer.sv"
	`include "Driver.sv"
	`include "Monitor.sv"
	`include "Subscriber.sv"
	`include "Scoreboard.sv"
	`include "Agent.sv"
	`include "Environment.sv"
	`include "Test.sv"

endpackage